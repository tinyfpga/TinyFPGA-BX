module TinyFPGA_B (
  output pin_pu,
  output pin_led
);
  assign pin_pu = 1'b0;
  assign pin_led = 1'b0;
endmodule
